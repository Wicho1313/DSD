module prioridad ( 
	num,
	cod
	) ;

input [8:0] num;
inout [3:0] cod;
