module conreg ( 
	clr,
	clk,
	e,
	c,
	q
	) ;

input  clr;
input  clk;
input [3:0] e;
input [2:0] c;
inout [3:0] q;
