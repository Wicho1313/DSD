module clock ( 
	t,
	clk,
	clr,
	pre,
	q,
	qn
	) ;

input  t;
input  clk;
input  clr;
input  pre;
inout  q;
inout  qn;
