module examen ( 
	clr,
	clk,
	c,
	q,
	disp
	) ;

input  clr;
input  clk;
input  c;
inout [2:0] q;
inout [6:0] disp;
