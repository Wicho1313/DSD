module contador ( 
	clk,
	clr,
	c,
	q
	) ;

input  clk;
input  clr;
input  c;
inout [7:0] q;
