module pseis ( 
	clr,
	clk,
	c,
	display
	) ;

input  clr;
input  clk;
input  c;
inout [6:0] display;
