--PRACTICA: 02_DSD
--AUTOR: 
--CODIGO: FF_SR

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFSR IS
PORT (
S,R,CLK,CLR,PRE: IN STD_LOGIC;
Q, NQ: INOUT STD_LOGIC
);
END FFSR;

ARCHITECTURE A_FFSR OF FFSR IS
SIGNAL AUX: STD_LOGIC;
BEGIN
AUX<=NOT(S OR (Q AND (NOT R)));
	PROCESS(S,R,CLK,CLR,PRE)
	BEGIN
		IF (CLR='0') THEN
			Q<='0';
			NQ<='1';
		ELSIF (CLK'EVENT AND CLK='1') THEN
			IF(PRE='1') THEN
				Q<='1';
				NQ<='0';
			ELSE 
				Q<= (S OR (Q AND (NOT R)));
				NQ<=((not q) or r)and (not s);
			END IF;
		END IF;
	END PROCESS;
END A_FFSR;