LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PRACTICA1 IS
PORT(
A,B,C,D,REF,SEL : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
DISPLAY: OUT STD_LOGIC_VECTOR (6 DOWNTO 0);
Z : INOUT  STD_LOGIC_VECTOR (1 DOWNTO 0));
END ENTITY;

--attribute pin_numbers of PRACTICA1: ENTITY IS
	--"A(1):1 A(0):2 B(1):3 B(0):4 C(1):5 C(0):6 D(1):7 D(0):8 SEL(1):9 SEL(0):10 REF(1):11 REF(0):14" 
--	& " DISPLAY(6):23 DISPLAY(5):22 DISPLAY(4):21 DISPLAY(3):20 DISPLAY(2):19 DISPLAY(1):18 DISPLAY(0):17 Z(1):16 Z(0):15";

--END PRACTICA1;


ARCHITECTURE A_PRAC1 OF PRACTICA1 IS 
	SIGNAL SAL: STD_LOGIC_VECTOR (2 DOWNTO 0);
	CONSTANT IGUAL: STD_LOGIC_VECTOR (6 DOWNTO 0):= "0111110";
	CONSTANT MAYOR: STD_LOGIC_VECTOR (6 DOWNTO 0):= "0011110";
	CONSTANT MENOR: STD_LOGIC_VECTOR (6 DOWNTO 0):= "0111100";

	BEGIN 


		PROCESS (SEL,A,B,C,D)
		BEGIN 
		CASE SEL IS 
		WHEN "00" => Z <= A;
		WHEN "01" => Z <= B;
		WHEN "10" => Z <= C;
		WHEN OTHERS => Z <= D;
		END CASE;
		END PROCESS;

		COMP: PROCESS (Z, REF)
		BEGIN
		IF(Z=REF) THEN 
			SAL <= "100";
		ELSIF( Z > REF) THEN 
			SAL <= "010";
		ELSE
			SAL <= "001";
			END IF;
		END PROCESS COMP ;


		DECO: PROCESS (SAL)
		BEGIN
		IF(SAL = "100") THEN 
			DISPLAY <= IGUAL;

		ELSIF (SAL = "010") THEN
			DISPLAY <= MAYOR; 

		ELSE 
			DISPLAY <= MENOR;
		END IF;

		END PROCESS DECO ; 
	END A_PRAC1;