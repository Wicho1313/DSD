module ffsr ( 
	s,
	r,
	clk,
	clr,
	pre,
	q,
	nq
	) ;

input  s;
input  r;
input  clk;
input  clr;
input  pre;
inout  q;
inout  nq;
